`define instr .lb(lb),.lbu(lbu),.lh(lh),.lhu(lhu),.lw(lw),.sb(sb),.sh(sh),.sw(sw),.add(add),.addu(addu),.subu(subu),.sub(sub),.mult(mult),.multu(multu),.div(div),.divu(divu),.sll(sll),.srl(srl),.sra(sra),.sllv(sllv),.srlv(srlv),.srav(srav),.And(And),.Or(Or),.Xor(Xor),.Nor(Nor),.addi(addi),.addiu(addiu),.andi(andi),.ori(ori),.xori(xori),.lui(lui),.slt(slt),.slti(slti),.sltiu(sltiu),.sltu(sltu),.beq(beq),.bne(bne),.blez(blez),.bgtz(bgtz),.bltz(bltz),.bgez(bgez),.j(j),.jal(jal),.jalr(jalr),.jr(jr),.mfhi(mfhi),.mflo(mflo),.mthi(mthi),.mtlo(mtlo),.eret(eret),.mtc0(mtc0),.mfc0(mfc0),.wrong(wrong)
`define rs 25:21
`define rt 20:16
`define rd 15:11
`define op 31:26
`define fuc 5:0