`define instr .addu(addu),.subu(subu),.lw(lw),.sw(sw),.beq(beq),.lui(lui),.jal(jal),.jr(jr),.ori(ori),.j(j),.cmco(cmco)
`define rs 25:21
`define rt 20:16
`define rd 15:11