`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   11:51:55 10/24/2020
// Design Name:   gray
// Module Name:   D:/verilog/gray/test.v
// Project Name:  gray
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: gray
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module test;

	// Inputs
	reg Clk;
	reg Reset;
	reg En;

	// Outputs
	wire [2:0] Output;
	wire Overflow;

	// Instantiate the Unit Under Test (UUT)
	gray uut (
		.Clk(Clk), 
		.Reset(Reset), 
		.En(En), 
		.Output(Output), 
		.Overflow(Overflow)
	);

	initial begin
		// Initialize Inputs
		Clk = 0;
		Reset = 0;
		En = 0;

		// Wait 100 ns for global reset to finish
		#100
      En =1;
      #10	
      En =1;
      #10
      En =1;
      #10
      En =1;
      #10		
		En =1;
      #10
		En =1;
      #10
		En =1;
      #10
		En =1;
      #10
		En =1;
      #10
		En =1;
      #10
		En =1;
		// Add stimulus here
end
     always #5 Clk = ~Clk;  
endmodule

