`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   10:18:42 09/19/2020
// Design Name:   cpu_checker
// Module Name:   D:/verilog/cpu/test2.v
// Project Name:  cpu
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: cpu_checker
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module test2;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	cpu_checker uut (
		.()
	);

	initial begin
		// Initialize Inputs
 
		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

